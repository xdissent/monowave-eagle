Double Balanced Multiplier
.CONTROL
run
.ENDC
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.SUBCKT OPAMP 1 2 101 102 81
.model NPN  NPN(BF=50000)
Q1 5 1 7 NPN
Q2 6 2 8 NPN
RC1 101 5 95.49
RC2 101 6 95.49
RE1 7 4 43.79
RE2 8 4 43.79
I1 4 102 0.001
G1 100 10 6 5 0.0104719
RP1 10 100 9.549MEG
CP1 10 100 0.0016667UF
EOUT 80 100 10 100 1
RO 80 81 100
RREF1 101 103 100K
RREF2 103 102 100K
EREF 100 0 103 0 1
R100 100 0 1MEG
.ENDS
CC1 MOD N$13 10uF
CC2 N$14 INVMOD 10uF
.TRAN 1uS 100mS
.CONTROL
plot OUT
.ENDC
Q1 COL1 N$3 N$1 2N3904
Q2 COL2 N$4 N$1 2N3904
Q3 COL1 N$5 N$2 2N3904
Q4 COL2 N$6 N$2 2N3904
Q5 N$1 N$13 N$8 2N3904
Q6 N$2 N$14 N$9 2N3904
RR1 COL2 VCC 750
RR2 COL1 VCC 750
RR3 IN N$3 47
RR4 N$4 0 47
RR5 0 N$5 47
RR6 N$6 IN 47
RR7 VEE N$8 680
RR8 VEE N$9 680
RR9 N$13 VCC 3k
RR10 VEE N$13 1k
RR11 N$14 VCC 3k
RR12 VEE N$14 1k
RR13 0 MOD 100k
RR14 0 INVMOD 100k
RR15 COL2 N$7 20k
RR16 N$7 OUT 20k
RR17 COL1 N$10 15k
RR18 0 N$10 15k
XU1 N$10 N$7 VCC VEE OUT OPAMP
VVSIN1 IN 0 AC 1 SIN(0 1V 440Hz)
VVSIN2 MOD INVMOD SIN(0 100mV 10Hz)
VCC VCC 0 DC 15V
VEE VEE 0 DC -15V
