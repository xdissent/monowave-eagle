Lead MV
.CONTROL
run
.ENDC
.SUBCKT 12AX7 A G K
Bca ca 0 V=45+V(A,K)+95.43*V(G,K)
Bre re 0 V=URAMP(V(A,K)/5)-URAMP(V(A,K)/5-1)
Baa A K I=V(re)*1.147E-6*(URAMP(V(ca))^1.5)
Bgg G K I=5E-6*(URAMP(V(G,K)+0.2)^1.5)
Cgk G K 1.6P
Cgp G A 1.7P
Cpk A K 0.46P
.ENDS
.SUBCKT 12AX7 A G K
Bca ca 0 V=45+V(A,K)+95.43*V(G,K)
Bre re 0 V=URAMP(V(A,K)/5)-URAMP(V(A,K)/5-1)
Baa A K I=V(re)*1.147E-6*(URAMP(V(ca))^1.5)
Bgg G K I=5E-6*(URAMP(V(G,K)+0.2)^1.5)
Cgk G K 1.6P
Cgp G A 1.7P
Cpk A K 0.46P
.ENDS
CC1 N$3 0 680nF
CC2 N$4 N$11 22nF
CC3 N$11 N$5 470pF
CC4 N$5 IN2 1nF
CC5 N$8 N$10 22nf
CC6 N$10 IN3 470pF
CC7 OUT ROUT 22nF
.TRAN 1us 100ms
.CONTROL
plot IN IN2 IN3 ROUT
.ENDC
RR1 0 IN 1Meg
RR2 IN N$1 68k
RR3 0 N$3 2.7k
RR4 N$4 VCC 100k
RR5 N$5 N$11 470k
RR6CW N$5 IN2 31065.001000
RR6CCW IN2 0 968935.001000
RR7 0 N$7 10k
RR8 N$8 VCC 100k
RR9 IN3 N$10 470k
RR10 0 IN3 470k
RR11 0 N$13 820
RR12 N$12 VDD 100k
RR13 0 OUT 100k
RR14 0 ROUT 1Meg
XVR1A N$8 IN2 N$7 12AX7
XVR1B N$4 N$1 N$3 12AX7
XVR2A N$12 IN3 N$13 12AX7
XVR2B VDD N$12 OUT 12AX7
VVSIN1 IN 0 AC 1 SIN(0 1V 666Hz)
VCC VCC 0 DC 250V
VDD VDD 0 DC 260V
