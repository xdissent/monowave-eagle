Op Amp Buffers
.CONTROL
run
.ENDC
.SUBCKT OPAMP 1 2 101 102 81
.model NPN  NPN(BF=50000)
Q1 5 1 7 NPN
Q2 6 2 8 NPN
RC1 101 5 95.49
RC2 101 6 95.49
RE1 7 4 43.79
RE2 8 4 43.79
I1 4 102 0.001
G1 100 10 6 5 0.0104719
RP1 10 100 9.549MEG
CP1 10 100 0.0016667UF
EOUT 80 100 10 100 1
RO 80 81 100
RREF1 101 103 100K
RREF2 103 102 100K
EREF 100 0 103 0 1
R100 100 0 1MEG
.ENDS
.TRAN 1uS 10mS
.CONTROL
plot OUT INVOUT
.ENDC
R1 IN N$1 100k
R2 N$1 INVOUT 100k
XU1A IN OUT VCC VEE OUT OPAMP
XU1B 0 N$1 VCC VEE INVOUT OPAMP
VVSIN1 IN 0 AC 1 SIN(0 1V 1kHz)
VCC VCC 0 DC 10V
VEE VEE 0 DC -10V
