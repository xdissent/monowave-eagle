Phase Inverter
.CONTROL
run
.ENDC
.SUBCKT 12AX7 A G K
Bca ca 0 V=45+V(A,K)+95.43*V(G,K)
Bre re 0 V=URAMP(V(A,K)/5)-URAMP(V(A,K)/5-1)
Baa A K I=V(re)*1.147E-6*(URAMP(V(ca))^1.5)
Bgg G K I=5E-6*(URAMP(V(G,K)+0.2)^1.5)
Cgk G K 1.6P
Cgp G A 1.7P
Cpk A K 0.46P
.ENDS
CC1 AFAMPIN VR1AG 50nF
CC2 VR1AA VR1BG 50nF
CC3 N$7 0 50uF
CC4 VR1BA PHASEINVOUT1 50nF
CC5 N$9 PHASEINVOUT2 50nF
.TRAN 1us 100ms
.CONTROL
plot AFAMPIN VR1BG PHASEINVOUT1 PHASEINVOUT2
.ENDC
.TRAN 1uS 100mS
.CONTROL
plot VR1BA VR1BK 
.ENDC
RR1 VR1AA VCC 1Meg
RR2 VR1BA VCC 270k
RR3 0 VR1AK 5.6k
RR4 N$9 VR1BK 5.1k
RR5 0 VR1AG 1Meg
RR6 N$9 VR1BG 1.2Meg
RR7 0 N$9 270k
RR8 N$7 VR1AK 270
RR9 0 PHASEINVOUT2 220k
RR10 0 PHASEINVOUT1 220k
XVR1A VR1AA VR1AG VR1AK 12AX7
XVR1B VR1AA VR1AG VR1AK 12AX7
VVSIN1 AFAMPIN 0 AC 1 SIN(0 0.00001V 1kHz)
VCC VCC 0 DC 340V
