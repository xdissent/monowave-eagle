Potentiometer Tapers
.CONTROL
run
.ENDC
.TRAN 1uS 10mS
.CONTROL
plot LINOUT LOGOUT REVLOGOUT
.ENDC
RR1CW IN LINOUT 50000.001000
RR1CCW LINOUT 0 50000.001000
RR2CW IN LOGOUT 88656.001000
RR2CCW LOGOUT 0 11344.001000
RR3CW IN REVLOGOUT 11344.001000
RR3CCW REVLOGOUT 0 88656.001000
VVSIN1 IN 0 AC 1 SIN(0 1V 1kHz)
