BJT Differential Amplifier
.CONTROL
run
.ENDC
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.TRAN 1uS 10mS
.CONTROL
plot INVOUT OUT
.ENDC
Q1 INVOUT IN N$3 2N3904
Q2 OUT 0 N$2 2N3904
R1 INVOUT VCC 75k
R2 OUT VCC 75k
R3 N$1 N$3 1k
R4 N$1 N$2 1k
R5 VEE N$1 75k
VVSIN1 IN 0 AC 1 SIN(0 100mV 1kHz)
VCC VCC 0 DC 15V
VEE VEE 0 DC -15V
