Voltage Controlled Oscillator
.CONTROL
run
.ENDC
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.model 2N3904 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+ Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+ Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.SUBCKT OPAMP 1 2 101 102 81
.model NPN  NPN(BF=50000)
Q1 5 1 7 NPN
Q2 6 2 8 NPN
RC1 101 5 95.49
RC2 101 6 95.49
RE1 7 4 43.79
RE2 8 4 43.79
I1 4 102 0.001
G1 100 10 6 5 0.0104719
RP1 10 100 9.549MEG
CP1 10 100 0.0016667UF
EOUT 80 100 10 100 1
RO 80 81 100
RREF1 101 103 100K
RREF2 103 102 100K
EREF 100 0 103 0 1
R100 100 0 1MEG
.ENDS
CC1 TRIANGLE N$1 0.01uF
.CONTROL
tran 1000uS 10S
setplot tran1
plot TRIANGLE SQUARE
.ENDC
Q1 N$9 N$8 0 2N3904
Q2 VCC SQUARE N$7 2N3904
RR1 IN N$1 100k
RR2 IN N$2 49.9k
RR3 0 N$2 49.9k
RR4 N$9 N$1 49.9k
RR5 0 N$5 100k
RR6 N$5 VCC 100k
RR7 N$5 SQUARE 100k
RR8 N$8 N$7 10k
RR9 0 N$7 47k
XU1A N$2 N$1 VCC 0 TRIANGLE OPAMP
XU1B N$5 TRIANGLE VCC 0 SQUARE OPAMP
VCC VCC 0 10V
VIN IN 0 9V
