Cascaded Tube Stages
.CONTROL
run
.ENDC
CC1 N$1 G2 20nF
CC2 N$5 OUT 100nF
.TRAN 1uS 100mS
.CONTROL
plot G1 G2 OUT
.ENDC
RR1 N$1 VCC 100k
RR2 IN G1 68k
RR3 0 G1 1Meg
RR4 0 N$3 1.5k
RR5 0 G2 1Meg
RR6 N$5 VCC 100k
RR7 0 N$6 1.5k
RR8 0 OUT 1Meg
TEST
VVSIN1 IN 0 AC 1 SIN(0 1V 1kHz)
VCC VCC 0 DC 300V
